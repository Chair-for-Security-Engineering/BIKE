
----------------------------------------------------------------------------------
-- COPYRIGHT (c) 2020 ALL RIGHT RESERVED
--
-- COMPANY:           Ruhr-University Bochum, Chair for Security Engineering
-- AUTHOR:            Jan Richter-Brockmann
--
-- CREATE DATE:       2020-05-27
-- LAST CHANGES:      2020-05-27
-- MODULE NAME:       BIKE_SQUARING_K4_GENERIC
--
-- REVISION:          1.00 - File was automatically created by a Sage script for r=12323 and d=32.
--
-- LICENCE:           Please look at licence.txt
-- USAGE INFORMATION: Please look at readme.txt. If licence.txt or readme.txt
--                    are missing or	if you have questions regarding the code
--                    please contact Tim Güneysu (tim.gueneysu@rub.de) and
--                    Jan Richter-Brockmann (jan.richter-brockmann@rub.de)
--
-- THIS CODE AND INFORMATION ARE PROVIDED "AS IS" WITHOUT WARRANTY OF ANY 
-- KIND, EITHER EXPRESSED OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE
-- IMPLIED WARRANTIES OF MERCHANTABILITY AND/OR FITNESS FOR A
-- PARTICULAR PURPOSE.
----------------------------------------------------------------------------------
  
-- IMPORTS
----------------------------------------------------------------------------------
LIBRARY IEEE;
    USE IEEE.STD_LOGIC_1164.ALL;
    USE IEEE.NUMERIC_STD.ALL;

LIBRARY UNISIM;
    USE UNISIM.vcomponents.ALL;
LIBRARY UNIMACRO;
    USE unimacro.Vcomponents.ALL;

LIBRARY work;
    USE work.BIKE_SETTINGS.ALL;



-- ENTITY
----------------------------------------------------------------------------------
ENTITY BIKE_SQUARING_K4_GENERIC IS
  PORT (  
    -- CONTROL PORTS ----------------
    CLK             : IN  STD_LOGIC; 	
    RESET           : IN  STD_LOGIC;
    ENABLE          : IN  STD_LOGIC;
    DONE            : OUT STD_LOGIC;
    -- INPUT POL -------------------
    REN_IN          : OUT STD_LOGIC;
    ADDR_IN         : OUT STD_LOGIC_VECTOR(LOG2(WORDS)-1 DOWNTO 0);
    DIN_IN          : IN  STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
    -- OUTPUT POL ------------------
    WEN_OUT         : OUT STD_LOGIC;
    ADDR_OUT        : OUT STD_LOGIC_VECTOR(LOG2(WORDS)-1 DOWNTO 0);
    DOUT_OUT        : OUT STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0)
  );
END BIKE_SQUARING_K4_GENERIC;



-- ARCHITECTURE
----------------------------------------------------------------------------------
ARCHITECTURE Behavioral OF BIKE_SQUARING_K4_GENERIC IS
  
    
    
-- SIGNALS
----------------------------------------------------------------------------------
-- COUNTER
SIGNAL CNT_RST                          : STD_LOGIC;
SIGNAL CNT_EN                           : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL CNT_OUT_0                        : STD_LOGIC_VECTOR(LOG2(WORDS)-1 DOWNTO 0);
SIGNAL CNT_OUT_1                        : STD_LOGIC_VECTOR(LOG2(WORDS)-1 DOWNTO 0);
SIGNAL CNT_OUT_2                        : STD_LOGIC_VECTOR(LOG2(WORDS)-1 DOWNTO 0);
SIGNAL CNT_OUT_3                        : STD_LOGIC_VECTOR(LOG2(WORDS)-1 DOWNTO 0);
SIGNAL CNT_OUT_4                        : STD_LOGIC_VECTOR(LOG2(WORDS)-1 DOWNTO 0);
SIGNAL CNT_OUT_5                        : STD_LOGIC_VECTOR(LOG2(WORDS)-1 DOWNTO 0);
SIGNAL CNT_OUT_6                        : STD_LOGIC_VECTOR(LOG2(WORDS)-1 DOWNTO 0);
SIGNAL CNT_OUT_7                        : STD_LOGIC_VECTOR(LOG2(WORDS)-1 DOWNTO 0);
SIGNAL CNT_OUT_8                        : STD_LOGIC_VECTOR(LOG2(WORDS)-1 DOWNTO 0);
SIGNAL CNT_OUT_9                        : STD_LOGIC_VECTOR(LOG2(WORDS)-1 DOWNTO 0);
SIGNAL CNT_OUT_10                        : STD_LOGIC_VECTOR(LOG2(WORDS)-1 DOWNTO 0);
SIGNAL CNT_OUT_11                        : STD_LOGIC_VECTOR(LOG2(WORDS)-1 DOWNTO 0);
SIGNAL CNT_OUT_12                        : STD_LOGIC_VECTOR(LOG2(WORDS)-1 DOWNTO 0);
SIGNAL CNT_OUT_13                        : STD_LOGIC_VECTOR(LOG2(WORDS)-1 DOWNTO 0);
SIGNAL CNT_OUT_14                        : STD_LOGIC_VECTOR(LOG2(WORDS)-1 DOWNTO 0);
SIGNAL CNT_OUT_15                        : STD_LOGIC_VECTOR(LOG2(WORDS)-1 DOWNTO 0);

SIGNAL CNT_EN_OUT, CNT_RST_OUT          : STD_LOGIC;
SIGNAL CNT_DONE_OUT                     : STD_LOGIC;
SIGNAL CNT_OUT_OUT                      : STD_LOGIC_VECTOR(LOG2(WORDS)-1 DOWNTO 0);

SIGNAL CNT_EN_INIT, CNT_RST_INIT        : STD_LOGIC;
SIGNAL CNT_DONE_INIT                    : STD_LOGIC;
SIGNAL CNT_OUT_INIT                     : STD_LOGIC_VECTOR(LOG2(16)-1 DOWNTO 0);

-- REGISTER
SIGNAL SEL_REG_EN                       : STD_LOGIC;
SIGNAL REG_EN                           : STD_LOGIC_VECTOR(16 DOWNTO 0);
SIGNAL REG_IN                           : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL REG0_OUT                         : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL REG1_OUT                         : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL REG2_OUT                         : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL REG3_OUT                         : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL REG4_OUT                         : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL REG5_OUT                         : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL REG6_OUT                         : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL REG7_OUT                         : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL REG8_OUT                         : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL REG9_OUT                         : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL REG10_OUT                         : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL REG11_OUT                         : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL REG12_OUT                         : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL REG13_OUT                         : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL REG14_OUT                         : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL REG15_OUT                         : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL REG16_OUT                         : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);

-- CONTROL MEMORY
SIGNAL SEL_ADDR_EN                      : STD_LOGIC;
SIGNAL SEL_ADDR                         : STD_LOGIC_VECTOR(15 DOWNTO 0);

-- OUTPUT
SIGNAL DOUT_OUT_PRE                     : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_0, DOUT_PART_0              : STD_LOGIC_VECTOR(B_WIDTH/16-1 DOWNTO 0);
SIGNAL DOUT_1, DOUT_PART_1              : STD_LOGIC_VECTOR(B_WIDTH/16-1 DOWNTO 0);
SIGNAL DOUT_2, DOUT_PART_2              : STD_LOGIC_VECTOR(B_WIDTH/16-1 DOWNTO 0);
SIGNAL DOUT_3, DOUT_PART_3              : STD_LOGIC_VECTOR(B_WIDTH/16-1 DOWNTO 0);
SIGNAL DOUT_4, DOUT_PART_4              : STD_LOGIC_VECTOR(B_WIDTH/16-1 DOWNTO 0);
SIGNAL DOUT_5, DOUT_PART_5              : STD_LOGIC_VECTOR(B_WIDTH/16-1 DOWNTO 0);
SIGNAL DOUT_6, DOUT_PART_6              : STD_LOGIC_VECTOR(B_WIDTH/16-1 DOWNTO 0);
SIGNAL DOUT_7, DOUT_PART_7              : STD_LOGIC_VECTOR(B_WIDTH/16-1 DOWNTO 0);
SIGNAL DOUT_8, DOUT_PART_8              : STD_LOGIC_VECTOR(B_WIDTH/16-1 DOWNTO 0);
SIGNAL DOUT_9, DOUT_PART_9              : STD_LOGIC_VECTOR(B_WIDTH/16-1 DOWNTO 0);
SIGNAL DOUT_10, DOUT_PART_10              : STD_LOGIC_VECTOR(B_WIDTH/16-1 DOWNTO 0);
SIGNAL DOUT_11, DOUT_PART_11              : STD_LOGIC_VECTOR(B_WIDTH/16-1 DOWNTO 0);
SIGNAL DOUT_12, DOUT_PART_12              : STD_LOGIC_VECTOR(B_WIDTH/16-1 DOWNTO 0);
SIGNAL DOUT_13, DOUT_PART_13              : STD_LOGIC_VECTOR(B_WIDTH/16-1 DOWNTO 0);
SIGNAL DOUT_14, DOUT_PART_14              : STD_LOGIC_VECTOR(B_WIDTH/16-1 DOWNTO 0);
SIGNAL DOUT_15, DOUT_PART_15              : STD_LOGIC_VECTOR(B_WIDTH/16-1 DOWNTO 0);

SIGNAL DOUT_REG_COMB0_0                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB1_0                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB0_1                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB1_1                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB0_2                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB1_2                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB0_3                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB1_3                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB0_4                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB1_4                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB0_5                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB1_5                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB0_6                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB1_6                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB0_7                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB1_7                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB0_8                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB1_8                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB0_9                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB1_9                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB0_10                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB1_10                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB0_11                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB1_11                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB0_12                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB1_12                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB0_13                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB1_13                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB0_14                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB1_14                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB0_15                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);
SIGNAL DOUT_REG_COMB1_15                 : STD_LOGIC_VECTOR(B_WIDTH-1 DOWNTO 0);

SIGNAL WRITE_LAST                       : STD_LOGIC;
SIGNAL SEL_REG_OUT                      : STD_LOGIC_VECTOR(16 DOWNTO 0);
  
    
    
-- STATES
----------------------------------------------------------------------------------
TYPE STATES IS (S_RESET, S_INIT0, S_INIT1, S_WRITE, S_DONE);
SIGNAL STATE : STATES := S_RESET;



-- BEHAVIORAL
----------------------------------------------------------------------------------
BEGIN
  
    -- COUNTER -------------------------------------------------------------------
    CNT_DONE_OUT <= '0' WHEN CNT_OUT_OUT < STD_LOGIC_VECTOR(TO_UNSIGNED(WORDS-2, LOG2(WORDS))) ELSE '1';
    WRITE_LAST <= '1' WHEN CNT_OUT_OUT = STD_LOGIC_VECTOR(TO_UNSIGNED(WORDS-1, LOG2(WORDS))) ELSE '0';
    
    CNT_OUT : ENTITY work.BIKE_COUNTER_INC_STOP GENERIC MAP(SIZE => LOG2(WORDS), MAX_VALUE => WORDS)
    PORT MAP(CLK => CLK, EN => CNT_EN_OUT, RST => CNT_RST_OUT, CNT_OUT => CNT_OUT_OUT);
    
    CNT_DONE_INIT <= '0' WHEN CNT_OUT_INIT < STD_LOGIC_VECTOR(TO_UNSIGNED(15, LOG2(16))) ELSE '1';
    CNT_INIT : ENTITY work.BIKE_COUNTER_INC_STOP GENERIC MAP(SIZE => LOG2(16), MAX_VALUE => 15)
    PORT MAP(CLK => CLK, EN => CNT_EN_INIT, RST => CNT_RST_INIT, CNT_OUT => CNT_OUT_INIT);
    
    CNT_EN <= SEL_ADDR;
    
    CNT0 : ENTITY work.BIKE_COUNTER_INC_INIT GENERIC MAP(SIZE => LOG2(WORDS), MAX_VALUE => 362, INITIAL => 336)
    PORT MAP(CLK => CLK, EN => CNT_EN(0), RST => CNT_RST, CNT_OUT => CNT_OUT_0);
    CNT1 : ENTITY work.BIKE_COUNTER_INC_INIT GENERIC MAP(SIZE => LOG2(WORDS), MAX_VALUE => 337, INITIAL => 312)
    PORT MAP(CLK => CLK, EN => CNT_EN(1), RST => CNT_RST, CNT_OUT => CNT_OUT_1);
    CNT2 : ENTITY work.BIKE_COUNTER_INC_INIT GENERIC MAP(SIZE => LOG2(WORDS), MAX_VALUE => 313, INITIAL => 288)
    PORT MAP(CLK => CLK, EN => CNT_EN(2), RST => CNT_RST, CNT_OUT => CNT_OUT_2);
    CNT3 : ENTITY work.BIKE_COUNTER_INC_INIT GENERIC MAP(SIZE => LOG2(WORDS), MAX_VALUE => 289, INITIAL => 264)
    PORT MAP(CLK => CLK, EN => CNT_EN(3), RST => CNT_RST, CNT_OUT => CNT_OUT_3);
    CNT4 : ENTITY work.BIKE_COUNTER_INC_INIT GENERIC MAP(SIZE => LOG2(WORDS), MAX_VALUE => 265, INITIAL => 240)
    PORT MAP(CLK => CLK, EN => CNT_EN(4), RST => CNT_RST, CNT_OUT => CNT_OUT_4);
    CNT5 : ENTITY work.BIKE_COUNTER_INC_INIT GENERIC MAP(SIZE => LOG2(WORDS), MAX_VALUE => 241, INITIAL => 216)
    PORT MAP(CLK => CLK, EN => CNT_EN(5), RST => CNT_RST, CNT_OUT => CNT_OUT_5);
    CNT6 : ENTITY work.BIKE_COUNTER_INC_INIT GENERIC MAP(SIZE => LOG2(WORDS), MAX_VALUE => 217, INITIAL => 192)
    PORT MAP(CLK => CLK, EN => CNT_EN(6), RST => CNT_RST, CNT_OUT => CNT_OUT_6);
    CNT7 : ENTITY work.BIKE_COUNTER_INC_INIT GENERIC MAP(SIZE => LOG2(WORDS), MAX_VALUE => 193, INITIAL => 168)
    PORT MAP(CLK => CLK, EN => CNT_EN(7), RST => CNT_RST, CNT_OUT => CNT_OUT_7);
    CNT8 : ENTITY work.BIKE_COUNTER_INC_INIT GENERIC MAP(SIZE => LOG2(WORDS), MAX_VALUE => 169, INITIAL => 144)
    PORT MAP(CLK => CLK, EN => CNT_EN(8), RST => CNT_RST, CNT_OUT => CNT_OUT_8);
    CNT9 : ENTITY work.BIKE_COUNTER_INC_INIT GENERIC MAP(SIZE => LOG2(WORDS), MAX_VALUE => 145, INITIAL => 120)
    PORT MAP(CLK => CLK, EN => CNT_EN(9), RST => CNT_RST, CNT_OUT => CNT_OUT_9);
    CNT10 : ENTITY work.BIKE_COUNTER_INC_INIT GENERIC MAP(SIZE => LOG2(WORDS), MAX_VALUE => 121, INITIAL => 96)
    PORT MAP(CLK => CLK, EN => CNT_EN(10), RST => CNT_RST, CNT_OUT => CNT_OUT_10);
    CNT11 : ENTITY work.BIKE_COUNTER_INC_INIT GENERIC MAP(SIZE => LOG2(WORDS), MAX_VALUE => 97, INITIAL => 72)
    PORT MAP(CLK => CLK, EN => CNT_EN(11), RST => CNT_RST, CNT_OUT => CNT_OUT_11);
    CNT12 : ENTITY work.BIKE_COUNTER_INC_INIT GENERIC MAP(SIZE => LOG2(WORDS), MAX_VALUE => 73, INITIAL => 48)
    PORT MAP(CLK => CLK, EN => CNT_EN(12), RST => CNT_RST, CNT_OUT => CNT_OUT_12);
    CNT13 : ENTITY work.BIKE_COUNTER_INC_INIT GENERIC MAP(SIZE => LOG2(WORDS), MAX_VALUE => 49, INITIAL => 24)
    PORT MAP(CLK => CLK, EN => CNT_EN(13), RST => CNT_RST, CNT_OUT => CNT_OUT_13);
    CNT14 : ENTITY work.BIKE_COUNTER_INC_INIT GENERIC MAP(SIZE => LOG2(WORDS), MAX_VALUE => 386, INITIAL => 361)
    PORT MAP(CLK => CLK, EN => CNT_EN(14), RST => CNT_RST, CNT_OUT => CNT_OUT_14);
    CNT15 : ENTITY work.BIKE_COUNTER_INC_INIT GENERIC MAP(SIZE => LOG2(WORDS), MAX_VALUE => 25, INITIAL => 0)
    PORT MAP(CLK => CLK, EN => CNT_EN(15), RST => CNT_RST, CNT_OUT => CNT_OUT_15);  
    ------------------------------------------------------------------------------


    -- OUTPUT --------------------------------------------------------------------
    ADDR_OUT <= CNT_OUT_OUT;
    
    -- special case for the polynomial's last msbs
    DOUT_OUT <= DOUT_OUT_PRE WHEN WRITE_LAST = '0' ELSE (B_WIDTH-1 DOWNTO OVERHANG => '0') & DOUT_OUT_PRE(OVERHANG-1 DOWNTO 0);
    
    -- spread output
    DOUT_ASSIGN : FOR I IN 0 TO B_WIDTH/16-1 GENERATE
      DOUT_OUT_PRE(16*I+0)   <= DOUT_0(I);
      DOUT_OUT_PRE(16*I+1)   <= DOUT_1(I);
      DOUT_OUT_PRE(16*I+2)   <= DOUT_2(I);
      DOUT_OUT_PRE(16*I+3)   <= DOUT_3(I);
      DOUT_OUT_PRE(16*I+4)   <= DOUT_4(I);
      DOUT_OUT_PRE(16*I+5)   <= DOUT_5(I);
      DOUT_OUT_PRE(16*I+6)   <= DOUT_6(I);
      DOUT_OUT_PRE(16*I+7)   <= DOUT_7(I);
      DOUT_OUT_PRE(16*I+8)   <= DOUT_8(I);
      DOUT_OUT_PRE(16*I+9)   <= DOUT_9(I);
      DOUT_OUT_PRE(16*I+10)   <= DOUT_10(I);
      DOUT_OUT_PRE(16*I+11)   <= DOUT_11(I);
      DOUT_OUT_PRE(16*I+12)   <= DOUT_12(I);
      DOUT_OUT_PRE(16*I+13)   <= DOUT_13(I);
      DOUT_OUT_PRE(16*I+14)   <= DOUT_14(I);
      DOUT_OUT_PRE(16*I+15)   <= DOUT_15(I);
    END GENERATE;

    
    -- assignment for DOUT_0
    DOUT_0 <= DOUT_PART_0;
    WITH SEL_ADDR SELECT DOUT_PART_0 <=
      DOUT_REG_COMB0_0(1*B_WIDTH/16-1+0 DOWNTO 0*B_WIDTH/16+0) WHEN "0000000000000010",
      DOUT_REG_COMB0_0(2*B_WIDTH/16-1+0 DOWNTO 1*B_WIDTH/16+0) WHEN "0000000000000100",
      DOUT_REG_COMB0_0(3*B_WIDTH/16-1+0 DOWNTO 2*B_WIDTH/16+0) WHEN "0000000000001000",
      DOUT_REG_COMB0_0(4*B_WIDTH/16-1+0 DOWNTO 3*B_WIDTH/16+0) WHEN "0000000000010000",
      DOUT_REG_COMB0_0(5*B_WIDTH/16-1+0 DOWNTO 4*B_WIDTH/16+0) WHEN "0000000000100000",
      DOUT_REG_COMB0_0(6*B_WIDTH/16-1+0 DOWNTO 5*B_WIDTH/16+0) WHEN "0000000001000000",
      DOUT_REG_COMB0_0(7*B_WIDTH/16-1+0 DOWNTO 6*B_WIDTH/16+0) WHEN "0000000010000000",
      DOUT_REG_COMB0_0(8*B_WIDTH/16-1+0 DOWNTO 7*B_WIDTH/16+0) WHEN "0000000100000000",
      DOUT_REG_COMB0_0(9*B_WIDTH/16-1+0 DOWNTO 8*B_WIDTH/16+0) WHEN "0000001000000000",
      DOUT_REG_COMB0_0(10*B_WIDTH/16-1+0 DOWNTO 9*B_WIDTH/16+0) WHEN "0000010000000000",
      DOUT_REG_COMB0_0(11*B_WIDTH/16-1+0 DOWNTO 10*B_WIDTH/16+0) WHEN "0000100000000000",
      DOUT_REG_COMB0_0(12*B_WIDTH/16-1+0 DOWNTO 11*B_WIDTH/16+0) WHEN "0001000000000000",
      DOUT_REG_COMB0_0(13*B_WIDTH/16-1+0 DOWNTO 12*B_WIDTH/16+0) WHEN "0010000000000000",
      DOUT_REG_COMB0_0(14*B_WIDTH/16-1+0 DOWNTO 13*B_WIDTH/16+0) WHEN "0100000000000000",
      DOUT_REG_COMB0_0(15*B_WIDTH/16-1+0 DOWNTO 14*B_WIDTH/16+0) WHEN "1000000000000000",
      DOUT_REG_COMB0_0(16*B_WIDTH/16-1+0 DOWNTO 15*B_WIDTH/16+0) WHEN "0000000000000001",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB0_0 <=
      REG15_OUT WHEN "00000000000000001",
      REG14_OUT WHEN "00000000000000010",
      REG13_OUT WHEN "00000000000000100",
      REG12_OUT WHEN "00000000000001000",
      REG11_OUT WHEN "00000000000010000",
      REG10_OUT WHEN "00000000000100000",
      REG9_OUT WHEN "00000000001000000",
      REG8_OUT WHEN "00000000010000000",
      REG7_OUT WHEN "00000000100000000",
      REG6_OUT WHEN "00000001000000000",
      REG5_OUT WHEN "00000010000000000",
      REG4_OUT WHEN "00000100000000000",
      REG3_OUT WHEN "00001000000000000",
      REG2_OUT WHEN "00010000000000000",
      REG1_OUT WHEN "00100000000000000",
      REG0_OUT WHEN "01000000000000000",
      REG16_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB1_0 <=
      REG14_OUT WHEN "00000000000000001",
      REG13_OUT WHEN "00000000000000010",
      REG12_OUT WHEN "00000000000000100",
      REG11_OUT WHEN "00000000000001000",
      REG10_OUT WHEN "00000000000010000",
      REG9_OUT WHEN "00000000000100000",
      REG8_OUT WHEN "00000000001000000",
      REG7_OUT WHEN "00000000010000000",
      REG6_OUT WHEN "00000000100000000",
      REG5_OUT WHEN "00000001000000000",
      REG4_OUT WHEN "00000010000000000",
      REG3_OUT WHEN "00000100000000000",
      REG2_OUT WHEN "00001000000000000",
      REG1_OUT WHEN "00010000000000000",
      REG0_OUT WHEN "00100000000000000",
      REG16_OUT WHEN "01000000000000000",
      REG15_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 



    -- assignment for DOUT_1
    DOUT_1 <= DOUT_PART_1;
    WITH SEL_ADDR SELECT DOUT_PART_1 <=
      DOUT_REG_COMB0_1(6*B_WIDTH/16-1+1 DOWNTO 5*B_WIDTH/16+1) WHEN "0000000000000010",
      DOUT_REG_COMB0_1(7*B_WIDTH/16-1+1 DOWNTO 6*B_WIDTH/16+1) WHEN "0000000000000100",
      DOUT_REG_COMB0_1(8*B_WIDTH/16-1+1 DOWNTO 7*B_WIDTH/16+1) WHEN "0000000000001000",
      DOUT_REG_COMB0_1(9*B_WIDTH/16-1+1 DOWNTO 8*B_WIDTH/16+1) WHEN "0000000000010000",
      DOUT_REG_COMB0_1(10*B_WIDTH/16-1+1 DOWNTO 9*B_WIDTH/16+1) WHEN "0000000000100000",
      DOUT_REG_COMB0_1(11*B_WIDTH/16-1+1 DOWNTO 10*B_WIDTH/16+1) WHEN "0000000001000000",
      DOUT_REG_COMB0_1(12*B_WIDTH/16-1+1 DOWNTO 11*B_WIDTH/16+1) WHEN "0000000010000000",
      DOUT_REG_COMB0_1(13*B_WIDTH/16-1+1 DOWNTO 12*B_WIDTH/16+1) WHEN "0000000100000000",
      DOUT_REG_COMB0_1(14*B_WIDTH/16-1+1 DOWNTO 13*B_WIDTH/16+1) WHEN "0000001000000000",
      DOUT_REG_COMB0_1(15*B_WIDTH/16-1+1 DOWNTO 14*B_WIDTH/16+1) WHEN "0000010000000000",
      DOUT_REG_COMB1_1(0 DOWNTO 0) & DOUT_REG_COMB0_1(31 DOWNTO 15*B_WIDTH/16+1) WHEN "0000100000000000",
      DOUT_REG_COMB1_1(1*B_WIDTH/16-1+1 DOWNTO 0*B_WIDTH/16+1) WHEN "0001000000000000",
      DOUT_REG_COMB1_1(2*B_WIDTH/16-1+1 DOWNTO 1*B_WIDTH/16+1) WHEN "0010000000000000",
      DOUT_REG_COMB1_1(3*B_WIDTH/16-1+1 DOWNTO 2*B_WIDTH/16+1) WHEN "0100000000000000",
      DOUT_REG_COMB1_1(4*B_WIDTH/16-1+1 DOWNTO 3*B_WIDTH/16+1) WHEN "1000000000000000",
      DOUT_REG_COMB1_1(5*B_WIDTH/16-1+1 DOWNTO 4*B_WIDTH/16+1) WHEN "0000000000000001",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB0_1 <=
      REG9_OUT WHEN "00000000000000001",
      REG8_OUT WHEN "00000000000000010",
      REG7_OUT WHEN "00000000000000100",
      REG6_OUT WHEN "00000000000001000",
      REG5_OUT WHEN "00000000000010000",
      REG4_OUT WHEN "00000000000100000",
      REG3_OUT WHEN "00000000001000000",
      REG2_OUT WHEN "00000000010000000",
      REG1_OUT WHEN "00000000100000000",
      REG0_OUT WHEN "00000001000000000",
      REG16_OUT WHEN "00000010000000000",
      REG15_OUT WHEN "00000100000000000",
      REG14_OUT WHEN "00001000000000000",
      REG13_OUT WHEN "00010000000000000",
      REG12_OUT WHEN "00100000000000000",
      REG11_OUT WHEN "01000000000000000",
      REG10_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB1_1 <=
      REG8_OUT WHEN "00000000000000001",
      REG7_OUT WHEN "00000000000000010",
      REG6_OUT WHEN "00000000000000100",
      REG5_OUT WHEN "00000000000001000",
      REG4_OUT WHEN "00000000000010000",
      REG3_OUT WHEN "00000000000100000",
      REG2_OUT WHEN "00000000001000000",
      REG1_OUT WHEN "00000000010000000",
      REG0_OUT WHEN "00000000100000000",
      REG16_OUT WHEN "00000001000000000",
      REG15_OUT WHEN "00000010000000000",
      REG14_OUT WHEN "00000100000000000",
      REG13_OUT WHEN "00001000000000000",
      REG12_OUT WHEN "00010000000000000",
      REG11_OUT WHEN "00100000000000000",
      REG10_OUT WHEN "01000000000000000",
      REG9_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 



    -- assignment for DOUT_2
    DOUT_2 <= DOUT_PART_2;
    WITH SEL_ADDR SELECT DOUT_PART_2 <=
      DOUT_REG_COMB0_2(12*B_WIDTH/16-1+0 DOWNTO 11*B_WIDTH/16+0) WHEN "0000000000000010",
      DOUT_REG_COMB0_2(13*B_WIDTH/16-1+0 DOWNTO 12*B_WIDTH/16+0) WHEN "0000000000000100",
      DOUT_REG_COMB0_2(14*B_WIDTH/16-1+0 DOWNTO 13*B_WIDTH/16+0) WHEN "0000000000001000",
      DOUT_REG_COMB0_2(15*B_WIDTH/16-1+0 DOWNTO 14*B_WIDTH/16+0) WHEN "0000000000010000",
      DOUT_REG_COMB0_2(16*B_WIDTH/16-1+0 DOWNTO 15*B_WIDTH/16+0) WHEN "0000000000100000",
      DOUT_REG_COMB1_2(1*B_WIDTH/16-1+0 DOWNTO 0*B_WIDTH/16+0) WHEN "0000000001000000",
      DOUT_REG_COMB1_2(2*B_WIDTH/16-1+0 DOWNTO 1*B_WIDTH/16+0) WHEN "0000000010000000",
      DOUT_REG_COMB1_2(3*B_WIDTH/16-1+0 DOWNTO 2*B_WIDTH/16+0) WHEN "0000000100000000",
      DOUT_REG_COMB1_2(4*B_WIDTH/16-1+0 DOWNTO 3*B_WIDTH/16+0) WHEN "0000001000000000",
      DOUT_REG_COMB1_2(5*B_WIDTH/16-1+0 DOWNTO 4*B_WIDTH/16+0) WHEN "0000010000000000",
      DOUT_REG_COMB1_2(6*B_WIDTH/16-1+0 DOWNTO 5*B_WIDTH/16+0) WHEN "0000100000000000",
      DOUT_REG_COMB1_2(7*B_WIDTH/16-1+0 DOWNTO 6*B_WIDTH/16+0) WHEN "0001000000000000",
      DOUT_REG_COMB1_2(8*B_WIDTH/16-1+0 DOWNTO 7*B_WIDTH/16+0) WHEN "0010000000000000",
      DOUT_REG_COMB1_2(9*B_WIDTH/16-1+0 DOWNTO 8*B_WIDTH/16+0) WHEN "0100000000000000",
      DOUT_REG_COMB1_2(10*B_WIDTH/16-1+0 DOWNTO 9*B_WIDTH/16+0) WHEN "1000000000000000",
      DOUT_REG_COMB1_2(11*B_WIDTH/16-1+0 DOWNTO 10*B_WIDTH/16+0) WHEN "0000000000000001",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB0_2 <=
      REG4_OUT WHEN "00000000000000001",
      REG3_OUT WHEN "00000000000000010",
      REG2_OUT WHEN "00000000000000100",
      REG1_OUT WHEN "00000000000001000",
      REG0_OUT WHEN "00000000000010000",
      REG16_OUT WHEN "00000000000100000",
      REG15_OUT WHEN "00000000001000000",
      REG14_OUT WHEN "00000000010000000",
      REG13_OUT WHEN "00000000100000000",
      REG12_OUT WHEN "00000001000000000",
      REG11_OUT WHEN "00000010000000000",
      REG10_OUT WHEN "00000100000000000",
      REG9_OUT WHEN "00001000000000000",
      REG8_OUT WHEN "00010000000000000",
      REG7_OUT WHEN "00100000000000000",
      REG6_OUT WHEN "01000000000000000",
      REG5_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB1_2 <=
      REG3_OUT WHEN "00000000000000001",
      REG2_OUT WHEN "00000000000000010",
      REG1_OUT WHEN "00000000000000100",
      REG0_OUT WHEN "00000000000001000",
      REG16_OUT WHEN "00000000000010000",
      REG15_OUT WHEN "00000000000100000",
      REG14_OUT WHEN "00000000001000000",
      REG13_OUT WHEN "00000000010000000",
      REG12_OUT WHEN "00000000100000000",
      REG11_OUT WHEN "00000001000000000",
      REG10_OUT WHEN "00000010000000000",
      REG9_OUT WHEN "00000100000000000",
      REG8_OUT WHEN "00001000000000000",
      REG7_OUT WHEN "00010000000000000",
      REG6_OUT WHEN "00100000000000000",
      REG5_OUT WHEN "01000000000000000",
      REG4_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 



    -- assignment for DOUT_3
    DOUT_3 <= DOUT_PART_3;
    WITH SEL_ADDR SELECT DOUT_PART_3 <=
      DOUT_REG_COMB0_3(1*B_WIDTH/16-1+1 DOWNTO 0*B_WIDTH/16+1) WHEN "0000000000000010",
      DOUT_REG_COMB0_3(2*B_WIDTH/16-1+1 DOWNTO 1*B_WIDTH/16+1) WHEN "0000000000000100",
      DOUT_REG_COMB0_3(3*B_WIDTH/16-1+1 DOWNTO 2*B_WIDTH/16+1) WHEN "0000000000001000",
      DOUT_REG_COMB0_3(4*B_WIDTH/16-1+1 DOWNTO 3*B_WIDTH/16+1) WHEN "0000000000010000",
      DOUT_REG_COMB0_3(5*B_WIDTH/16-1+1 DOWNTO 4*B_WIDTH/16+1) WHEN "0000000000100000",
      DOUT_REG_COMB0_3(6*B_WIDTH/16-1+1 DOWNTO 5*B_WIDTH/16+1) WHEN "0000000001000000",
      DOUT_REG_COMB0_3(7*B_WIDTH/16-1+1 DOWNTO 6*B_WIDTH/16+1) WHEN "0000000010000000",
      DOUT_REG_COMB0_3(8*B_WIDTH/16-1+1 DOWNTO 7*B_WIDTH/16+1) WHEN "0000000100000000",
      DOUT_REG_COMB0_3(9*B_WIDTH/16-1+1 DOWNTO 8*B_WIDTH/16+1) WHEN "0000001000000000",
      DOUT_REG_COMB0_3(10*B_WIDTH/16-1+1 DOWNTO 9*B_WIDTH/16+1) WHEN "0000010000000000",
      DOUT_REG_COMB0_3(11*B_WIDTH/16-1+1 DOWNTO 10*B_WIDTH/16+1) WHEN "0000100000000000",
      DOUT_REG_COMB0_3(12*B_WIDTH/16-1+1 DOWNTO 11*B_WIDTH/16+1) WHEN "0001000000000000",
      DOUT_REG_COMB0_3(13*B_WIDTH/16-1+1 DOWNTO 12*B_WIDTH/16+1) WHEN "0010000000000000",
      DOUT_REG_COMB0_3(14*B_WIDTH/16-1+1 DOWNTO 13*B_WIDTH/16+1) WHEN "0100000000000000",
      DOUT_REG_COMB0_3(15*B_WIDTH/16-1+1 DOWNTO 14*B_WIDTH/16+1) WHEN "1000000000000000",
      DOUT_REG_COMB1_3(0 DOWNTO 0) & DOUT_REG_COMB0_3(31 DOWNTO 15*B_WIDTH/16+1) WHEN "0000000000000001",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB0_3 <=
      REG14_OUT WHEN "00000000000000001",
      REG13_OUT WHEN "00000000000000010",
      REG12_OUT WHEN "00000000000000100",
      REG11_OUT WHEN "00000000000001000",
      REG10_OUT WHEN "00000000000010000",
      REG9_OUT WHEN "00000000000100000",
      REG8_OUT WHEN "00000000001000000",
      REG7_OUT WHEN "00000000010000000",
      REG6_OUT WHEN "00000000100000000",
      REG5_OUT WHEN "00000001000000000",
      REG4_OUT WHEN "00000010000000000",
      REG3_OUT WHEN "00000100000000000",
      REG2_OUT WHEN "00001000000000000",
      REG1_OUT WHEN "00010000000000000",
      REG0_OUT WHEN "00100000000000000",
      REG16_OUT WHEN "01000000000000000",
      REG15_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB1_3 <=
      REG13_OUT WHEN "00000000000000001",
      REG12_OUT WHEN "00000000000000010",
      REG11_OUT WHEN "00000000000000100",
      REG10_OUT WHEN "00000000000001000",
      REG9_OUT WHEN "00000000000010000",
      REG8_OUT WHEN "00000000000100000",
      REG7_OUT WHEN "00000000001000000",
      REG6_OUT WHEN "00000000010000000",
      REG5_OUT WHEN "00000000100000000",
      REG4_OUT WHEN "00000001000000000",
      REG3_OUT WHEN "00000010000000000",
      REG2_OUT WHEN "00000100000000000",
      REG1_OUT WHEN "00001000000000000",
      REG0_OUT WHEN "00010000000000000",
      REG16_OUT WHEN "00100000000000000",
      REG15_OUT WHEN "01000000000000000",
      REG14_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 



    -- assignment for DOUT_4
    DOUT_4 <= DOUT_PART_4;
    WITH SEL_ADDR SELECT DOUT_PART_4 <=
      DOUT_REG_COMB0_4(5*B_WIDTH/16-1+1 DOWNTO 4*B_WIDTH/16+1) WHEN "0000000000000010",
      DOUT_REG_COMB0_4(6*B_WIDTH/16-1+1 DOWNTO 5*B_WIDTH/16+1) WHEN "0000000000000100",
      DOUT_REG_COMB0_4(7*B_WIDTH/16-1+1 DOWNTO 6*B_WIDTH/16+1) WHEN "0000000000001000",
      DOUT_REG_COMB0_4(8*B_WIDTH/16-1+1 DOWNTO 7*B_WIDTH/16+1) WHEN "0000000000010000",
      DOUT_REG_COMB0_4(9*B_WIDTH/16-1+1 DOWNTO 8*B_WIDTH/16+1) WHEN "0000000000100000",
      DOUT_REG_COMB0_4(10*B_WIDTH/16-1+1 DOWNTO 9*B_WIDTH/16+1) WHEN "0000000001000000",
      DOUT_REG_COMB0_4(11*B_WIDTH/16-1+1 DOWNTO 10*B_WIDTH/16+1) WHEN "0000000010000000",
      DOUT_REG_COMB0_4(12*B_WIDTH/16-1+1 DOWNTO 11*B_WIDTH/16+1) WHEN "0000000100000000",
      DOUT_REG_COMB0_4(13*B_WIDTH/16-1+1 DOWNTO 12*B_WIDTH/16+1) WHEN "0000001000000000",
      DOUT_REG_COMB0_4(14*B_WIDTH/16-1+1 DOWNTO 13*B_WIDTH/16+1) WHEN "0000010000000000",
      DOUT_REG_COMB0_4(15*B_WIDTH/16-1+1 DOWNTO 14*B_WIDTH/16+1) WHEN "0000100000000000",
      DOUT_REG_COMB1_4(0 DOWNTO 0) & DOUT_REG_COMB0_4(31 DOWNTO 15*B_WIDTH/16+1) WHEN "0001000000000000",
      DOUT_REG_COMB1_4(1*B_WIDTH/16-1+1 DOWNTO 0*B_WIDTH/16+1) WHEN "0010000000000000",
      DOUT_REG_COMB1_4(2*B_WIDTH/16-1+1 DOWNTO 1*B_WIDTH/16+1) WHEN "0100000000000000",
      DOUT_REG_COMB1_4(3*B_WIDTH/16-1+1 DOWNTO 2*B_WIDTH/16+1) WHEN "1000000000000000",
      DOUT_REG_COMB1_4(4*B_WIDTH/16-1+1 DOWNTO 3*B_WIDTH/16+1) WHEN "0000000000000001",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB0_4 <=
      REG10_OUT WHEN "00000000000000001",
      REG9_OUT WHEN "00000000000000010",
      REG8_OUT WHEN "00000000000000100",
      REG7_OUT WHEN "00000000000001000",
      REG6_OUT WHEN "00000000000010000",
      REG5_OUT WHEN "00000000000100000",
      REG4_OUT WHEN "00000000001000000",
      REG3_OUT WHEN "00000000010000000",
      REG2_OUT WHEN "00000000100000000",
      REG1_OUT WHEN "00000001000000000",
      REG0_OUT WHEN "00000010000000000",
      REG16_OUT WHEN "00000100000000000",
      REG15_OUT WHEN "00001000000000000",
      REG14_OUT WHEN "00010000000000000",
      REG13_OUT WHEN "00100000000000000",
      REG12_OUT WHEN "01000000000000000",
      REG11_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB1_4 <=
      REG9_OUT WHEN "00000000000000001",
      REG8_OUT WHEN "00000000000000010",
      REG7_OUT WHEN "00000000000000100",
      REG6_OUT WHEN "00000000000001000",
      REG5_OUT WHEN "00000000000010000",
      REG4_OUT WHEN "00000000000100000",
      REG3_OUT WHEN "00000000001000000",
      REG2_OUT WHEN "00000000010000000",
      REG1_OUT WHEN "00000000100000000",
      REG0_OUT WHEN "00000001000000000",
      REG16_OUT WHEN "00000010000000000",
      REG15_OUT WHEN "00000100000000000",
      REG14_OUT WHEN "00001000000000000",
      REG13_OUT WHEN "00010000000000000",
      REG12_OUT WHEN "00100000000000000",
      REG11_OUT WHEN "01000000000000000",
      REG10_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 



    -- assignment for DOUT_5
    DOUT_5 <= DOUT_PART_5;
    WITH SEL_ADDR SELECT DOUT_PART_5 <=
      DOUT_REG_COMB0_5(11*B_WIDTH/16-1+0 DOWNTO 10*B_WIDTH/16+0) WHEN "0000000000000010",
      DOUT_REG_COMB0_5(12*B_WIDTH/16-1+0 DOWNTO 11*B_WIDTH/16+0) WHEN "0000000000000100",
      DOUT_REG_COMB0_5(13*B_WIDTH/16-1+0 DOWNTO 12*B_WIDTH/16+0) WHEN "0000000000001000",
      DOUT_REG_COMB0_5(14*B_WIDTH/16-1+0 DOWNTO 13*B_WIDTH/16+0) WHEN "0000000000010000",
      DOUT_REG_COMB0_5(15*B_WIDTH/16-1+0 DOWNTO 14*B_WIDTH/16+0) WHEN "0000000000100000",
      DOUT_REG_COMB0_5(16*B_WIDTH/16-1+0 DOWNTO 15*B_WIDTH/16+0) WHEN "0000000001000000",
      DOUT_REG_COMB1_5(1*B_WIDTH/16-1+0 DOWNTO 0*B_WIDTH/16+0) WHEN "0000000010000000",
      DOUT_REG_COMB1_5(2*B_WIDTH/16-1+0 DOWNTO 1*B_WIDTH/16+0) WHEN "0000000100000000",
      DOUT_REG_COMB1_5(3*B_WIDTH/16-1+0 DOWNTO 2*B_WIDTH/16+0) WHEN "0000001000000000",
      DOUT_REG_COMB1_5(4*B_WIDTH/16-1+0 DOWNTO 3*B_WIDTH/16+0) WHEN "0000010000000000",
      DOUT_REG_COMB1_5(5*B_WIDTH/16-1+0 DOWNTO 4*B_WIDTH/16+0) WHEN "0000100000000000",
      DOUT_REG_COMB1_5(6*B_WIDTH/16-1+0 DOWNTO 5*B_WIDTH/16+0) WHEN "0001000000000000",
      DOUT_REG_COMB1_5(7*B_WIDTH/16-1+0 DOWNTO 6*B_WIDTH/16+0) WHEN "0010000000000000",
      DOUT_REG_COMB1_5(8*B_WIDTH/16-1+0 DOWNTO 7*B_WIDTH/16+0) WHEN "0100000000000000",
      DOUT_REG_COMB1_5(9*B_WIDTH/16-1+0 DOWNTO 8*B_WIDTH/16+0) WHEN "1000000000000000",
      DOUT_REG_COMB1_5(10*B_WIDTH/16-1+0 DOWNTO 9*B_WIDTH/16+0) WHEN "0000000000000001",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB0_5 <=
      REG5_OUT WHEN "00000000000000001",
      REG4_OUT WHEN "00000000000000010",
      REG3_OUT WHEN "00000000000000100",
      REG2_OUT WHEN "00000000000001000",
      REG1_OUT WHEN "00000000000010000",
      REG0_OUT WHEN "00000000000100000",
      REG16_OUT WHEN "00000000001000000",
      REG15_OUT WHEN "00000000010000000",
      REG14_OUT WHEN "00000000100000000",
      REG13_OUT WHEN "00000001000000000",
      REG12_OUT WHEN "00000010000000000",
      REG11_OUT WHEN "00000100000000000",
      REG10_OUT WHEN "00001000000000000",
      REG9_OUT WHEN "00010000000000000",
      REG8_OUT WHEN "00100000000000000",
      REG7_OUT WHEN "01000000000000000",
      REG6_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB1_5 <=
      REG4_OUT WHEN "00000000000000001",
      REG3_OUT WHEN "00000000000000010",
      REG2_OUT WHEN "00000000000000100",
      REG1_OUT WHEN "00000000000001000",
      REG0_OUT WHEN "00000000000010000",
      REG16_OUT WHEN "00000000000100000",
      REG15_OUT WHEN "00000000001000000",
      REG14_OUT WHEN "00000000010000000",
      REG13_OUT WHEN "00000000100000000",
      REG12_OUT WHEN "00000001000000000",
      REG11_OUT WHEN "00000010000000000",
      REG10_OUT WHEN "00000100000000000",
      REG9_OUT WHEN "00001000000000000",
      REG8_OUT WHEN "00010000000000000",
      REG7_OUT WHEN "00100000000000000",
      REG6_OUT WHEN "01000000000000000",
      REG5_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 



    -- assignment for DOUT_6
    DOUT_6 <= DOUT_PART_6;
    WITH SEL_ADDR SELECT DOUT_PART_6 <=
      DIN_IN(0 DOWNTO 0) & DOUT_REG_COMB0_6(31 DOWNTO 15*B_WIDTH/16+1) WHEN "0000000000000010",
      DOUT_REG_COMB1_6(1*B_WIDTH/16-1+1 DOWNTO 0*B_WIDTH/16+1) WHEN "0000000000000100",
      DOUT_REG_COMB1_6(2*B_WIDTH/16-1+1 DOWNTO 1*B_WIDTH/16+1) WHEN "0000000000001000",
      DOUT_REG_COMB1_6(3*B_WIDTH/16-1+1 DOWNTO 2*B_WIDTH/16+1) WHEN "0000000000010000",
      DOUT_REG_COMB1_6(4*B_WIDTH/16-1+1 DOWNTO 3*B_WIDTH/16+1) WHEN "0000000000100000",
      DOUT_REG_COMB1_6(5*B_WIDTH/16-1+1 DOWNTO 4*B_WIDTH/16+1) WHEN "0000000001000000",
      DOUT_REG_COMB1_6(6*B_WIDTH/16-1+1 DOWNTO 5*B_WIDTH/16+1) WHEN "0000000010000000",
      DOUT_REG_COMB1_6(7*B_WIDTH/16-1+1 DOWNTO 6*B_WIDTH/16+1) WHEN "0000000100000000",
      DOUT_REG_COMB1_6(8*B_WIDTH/16-1+1 DOWNTO 7*B_WIDTH/16+1) WHEN "0000001000000000",
      DOUT_REG_COMB1_6(9*B_WIDTH/16-1+1 DOWNTO 8*B_WIDTH/16+1) WHEN "0000010000000000",
      DOUT_REG_COMB1_6(10*B_WIDTH/16-1+1 DOWNTO 9*B_WIDTH/16+1) WHEN "0000100000000000",
      DOUT_REG_COMB1_6(11*B_WIDTH/16-1+1 DOWNTO 10*B_WIDTH/16+1) WHEN "0001000000000000",
      DOUT_REG_COMB1_6(12*B_WIDTH/16-1+1 DOWNTO 11*B_WIDTH/16+1) WHEN "0010000000000000",
      DOUT_REG_COMB1_6(13*B_WIDTH/16-1+1 DOWNTO 12*B_WIDTH/16+1) WHEN "0100000000000000",
      DOUT_REG_COMB1_6(14*B_WIDTH/16-1+1 DOWNTO 13*B_WIDTH/16+1) WHEN "1000000000000000",
      DOUT_REG_COMB1_6(15*B_WIDTH/16-1+1 DOWNTO 14*B_WIDTH/16+1) WHEN "0000000000000001",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB0_6 <=
      REG0_OUT WHEN "00000000000000001",
      REG16_OUT WHEN "00000000000000010",
      REG15_OUT WHEN "00000000000000100",
      REG14_OUT WHEN "00000000000001000",
      REG13_OUT WHEN "00000000000010000",
      REG12_OUT WHEN "00000000000100000",
      REG11_OUT WHEN "00000000001000000",
      REG10_OUT WHEN "00000000010000000",
      REG9_OUT WHEN "00000000100000000",
      REG8_OUT WHEN "00000001000000000",
      REG7_OUT WHEN "00000010000000000",
      REG6_OUT WHEN "00000100000000000",
      REG5_OUT WHEN "00001000000000000",
      REG4_OUT WHEN "00010000000000000",
      REG3_OUT WHEN "00100000000000000",
      REG2_OUT WHEN "01000000000000000",
      REG1_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB1_6 <=
      REG16_OUT WHEN "00000000000000001",
      REG15_OUT WHEN "00000000000000010",
      REG14_OUT WHEN "00000000000000100",
      REG13_OUT WHEN "00000000000001000",
      REG12_OUT WHEN "00000000000010000",
      REG11_OUT WHEN "00000000000100000",
      REG10_OUT WHEN "00000000001000000",
      REG9_OUT WHEN "00000000010000000",
      REG8_OUT WHEN "00000000100000000",
      REG7_OUT WHEN "00000001000000000",
      REG6_OUT WHEN "00000010000000000",
      REG5_OUT WHEN "00000100000000000",
      REG4_OUT WHEN "00001000000000000",
      REG3_OUT WHEN "00010000000000000",
      REG2_OUT WHEN "00100000000000000",
      REG1_OUT WHEN "01000000000000000",
      REG0_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 



    -- assignment for DOUT_7
    DOUT_7 <= DOUT_PART_7;
    WITH SEL_ADDR SELECT DOUT_PART_7 <=
      DOUT_REG_COMB0_7(4*B_WIDTH/16-1+1 DOWNTO 3*B_WIDTH/16+1) WHEN "0000000000000010",
      DOUT_REG_COMB0_7(5*B_WIDTH/16-1+1 DOWNTO 4*B_WIDTH/16+1) WHEN "0000000000000100",
      DOUT_REG_COMB0_7(6*B_WIDTH/16-1+1 DOWNTO 5*B_WIDTH/16+1) WHEN "0000000000001000",
      DOUT_REG_COMB0_7(7*B_WIDTH/16-1+1 DOWNTO 6*B_WIDTH/16+1) WHEN "0000000000010000",
      DOUT_REG_COMB0_7(8*B_WIDTH/16-1+1 DOWNTO 7*B_WIDTH/16+1) WHEN "0000000000100000",
      DOUT_REG_COMB0_7(9*B_WIDTH/16-1+1 DOWNTO 8*B_WIDTH/16+1) WHEN "0000000001000000",
      DOUT_REG_COMB0_7(10*B_WIDTH/16-1+1 DOWNTO 9*B_WIDTH/16+1) WHEN "0000000010000000",
      DOUT_REG_COMB0_7(11*B_WIDTH/16-1+1 DOWNTO 10*B_WIDTH/16+1) WHEN "0000000100000000",
      DOUT_REG_COMB0_7(12*B_WIDTH/16-1+1 DOWNTO 11*B_WIDTH/16+1) WHEN "0000001000000000",
      DOUT_REG_COMB0_7(13*B_WIDTH/16-1+1 DOWNTO 12*B_WIDTH/16+1) WHEN "0000010000000000",
      DOUT_REG_COMB0_7(14*B_WIDTH/16-1+1 DOWNTO 13*B_WIDTH/16+1) WHEN "0000100000000000",
      DOUT_REG_COMB0_7(15*B_WIDTH/16-1+1 DOWNTO 14*B_WIDTH/16+1) WHEN "0001000000000000",
      DOUT_REG_COMB1_7(0 DOWNTO 0) & DOUT_REG_COMB0_7(31 DOWNTO 15*B_WIDTH/16+1) WHEN "0010000000000000",
      DOUT_REG_COMB1_7(1*B_WIDTH/16-1+1 DOWNTO 0*B_WIDTH/16+1) WHEN "0100000000000000",
      DOUT_REG_COMB1_7(2*B_WIDTH/16-1+1 DOWNTO 1*B_WIDTH/16+1) WHEN "1000000000000000",
      DOUT_REG_COMB1_7(3*B_WIDTH/16-1+1 DOWNTO 2*B_WIDTH/16+1) WHEN "0000000000000001",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB0_7 <=
      REG11_OUT WHEN "00000000000000001",
      REG10_OUT WHEN "00000000000000010",
      REG9_OUT WHEN "00000000000000100",
      REG8_OUT WHEN "00000000000001000",
      REG7_OUT WHEN "00000000000010000",
      REG6_OUT WHEN "00000000000100000",
      REG5_OUT WHEN "00000000001000000",
      REG4_OUT WHEN "00000000010000000",
      REG3_OUT WHEN "00000000100000000",
      REG2_OUT WHEN "00000001000000000",
      REG1_OUT WHEN "00000010000000000",
      REG0_OUT WHEN "00000100000000000",
      REG16_OUT WHEN "00001000000000000",
      REG15_OUT WHEN "00010000000000000",
      REG14_OUT WHEN "00100000000000000",
      REG13_OUT WHEN "01000000000000000",
      REG12_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB1_7 <=
      REG10_OUT WHEN "00000000000000001",
      REG9_OUT WHEN "00000000000000010",
      REG8_OUT WHEN "00000000000000100",
      REG7_OUT WHEN "00000000000001000",
      REG6_OUT WHEN "00000000000010000",
      REG5_OUT WHEN "00000000000100000",
      REG4_OUT WHEN "00000000001000000",
      REG3_OUT WHEN "00000000010000000",
      REG2_OUT WHEN "00000000100000000",
      REG1_OUT WHEN "00000001000000000",
      REG0_OUT WHEN "00000010000000000",
      REG16_OUT WHEN "00000100000000000",
      REG15_OUT WHEN "00001000000000000",
      REG14_OUT WHEN "00010000000000000",
      REG13_OUT WHEN "00100000000000000",
      REG12_OUT WHEN "01000000000000000",
      REG11_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 



    -- assignment for DOUT_8
    DOUT_8 <= DOUT_PART_8;
    WITH SEL_ADDR SELECT DOUT_PART_8 <=
      DOUT_REG_COMB0_8(10*B_WIDTH/16-1+0 DOWNTO 9*B_WIDTH/16+0) WHEN "0000000000000010",
      DOUT_REG_COMB0_8(11*B_WIDTH/16-1+0 DOWNTO 10*B_WIDTH/16+0) WHEN "0000000000000100",
      DOUT_REG_COMB0_8(12*B_WIDTH/16-1+0 DOWNTO 11*B_WIDTH/16+0) WHEN "0000000000001000",
      DOUT_REG_COMB0_8(13*B_WIDTH/16-1+0 DOWNTO 12*B_WIDTH/16+0) WHEN "0000000000010000",
      DOUT_REG_COMB0_8(14*B_WIDTH/16-1+0 DOWNTO 13*B_WIDTH/16+0) WHEN "0000000000100000",
      DOUT_REG_COMB0_8(15*B_WIDTH/16-1+0 DOWNTO 14*B_WIDTH/16+0) WHEN "0000000001000000",
      DOUT_REG_COMB0_8(16*B_WIDTH/16-1+0 DOWNTO 15*B_WIDTH/16+0) WHEN "0000000010000000",
      DOUT_REG_COMB1_8(1*B_WIDTH/16-1+0 DOWNTO 0*B_WIDTH/16+0) WHEN "0000000100000000",
      DOUT_REG_COMB1_8(2*B_WIDTH/16-1+0 DOWNTO 1*B_WIDTH/16+0) WHEN "0000001000000000",
      DOUT_REG_COMB1_8(3*B_WIDTH/16-1+0 DOWNTO 2*B_WIDTH/16+0) WHEN "0000010000000000",
      DOUT_REG_COMB1_8(4*B_WIDTH/16-1+0 DOWNTO 3*B_WIDTH/16+0) WHEN "0000100000000000",
      DOUT_REG_COMB1_8(5*B_WIDTH/16-1+0 DOWNTO 4*B_WIDTH/16+0) WHEN "0001000000000000",
      DOUT_REG_COMB1_8(6*B_WIDTH/16-1+0 DOWNTO 5*B_WIDTH/16+0) WHEN "0010000000000000",
      DOUT_REG_COMB1_8(7*B_WIDTH/16-1+0 DOWNTO 6*B_WIDTH/16+0) WHEN "0100000000000000",
      DOUT_REG_COMB1_8(8*B_WIDTH/16-1+0 DOWNTO 7*B_WIDTH/16+0) WHEN "1000000000000000",
      DOUT_REG_COMB1_8(9*B_WIDTH/16-1+0 DOWNTO 8*B_WIDTH/16+0) WHEN "0000000000000001",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB0_8 <=
      REG6_OUT WHEN "00000000000000001",
      REG5_OUT WHEN "00000000000000010",
      REG4_OUT WHEN "00000000000000100",
      REG3_OUT WHEN "00000000000001000",
      REG2_OUT WHEN "00000000000010000",
      REG1_OUT WHEN "00000000000100000",
      REG0_OUT WHEN "00000000001000000",
      REG16_OUT WHEN "00000000010000000",
      REG15_OUT WHEN "00000000100000000",
      REG14_OUT WHEN "00000001000000000",
      REG13_OUT WHEN "00000010000000000",
      REG12_OUT WHEN "00000100000000000",
      REG11_OUT WHEN "00001000000000000",
      REG10_OUT WHEN "00010000000000000",
      REG9_OUT WHEN "00100000000000000",
      REG8_OUT WHEN "01000000000000000",
      REG7_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB1_8 <=
      REG5_OUT WHEN "00000000000000001",
      REG4_OUT WHEN "00000000000000010",
      REG3_OUT WHEN "00000000000000100",
      REG2_OUT WHEN "00000000000001000",
      REG1_OUT WHEN "00000000000010000",
      REG0_OUT WHEN "00000000000100000",
      REG16_OUT WHEN "00000000001000000",
      REG15_OUT WHEN "00000000010000000",
      REG14_OUT WHEN "00000000100000000",
      REG13_OUT WHEN "00000001000000000",
      REG12_OUT WHEN "00000010000000000",
      REG11_OUT WHEN "00000100000000000",
      REG10_OUT WHEN "00001000000000000",
      REG9_OUT WHEN "00010000000000000",
      REG8_OUT WHEN "00100000000000000",
      REG7_OUT WHEN "01000000000000000",
      REG6_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 



    -- assignment for DOUT_9
    DOUT_9 <= DOUT_PART_9;
    WITH SEL_ADDR SELECT DOUT_PART_9 <=
      DOUT_REG_COMB0_9(15*B_WIDTH/16-1+1 DOWNTO 14*B_WIDTH/16+1) WHEN "0000000000000010",
      DIN_IN(0 DOWNTO 0) & DOUT_REG_COMB0_9(31 DOWNTO 15*B_WIDTH/16+1) WHEN "0000000000000100",
      DOUT_REG_COMB1_9(1*B_WIDTH/16-1+1 DOWNTO 0*B_WIDTH/16+1) WHEN "0000000000001000",
      DOUT_REG_COMB1_9(2*B_WIDTH/16-1+1 DOWNTO 1*B_WIDTH/16+1) WHEN "0000000000010000",
      DOUT_REG_COMB1_9(3*B_WIDTH/16-1+1 DOWNTO 2*B_WIDTH/16+1) WHEN "0000000000100000",
      DOUT_REG_COMB1_9(4*B_WIDTH/16-1+1 DOWNTO 3*B_WIDTH/16+1) WHEN "0000000001000000",
      DOUT_REG_COMB1_9(5*B_WIDTH/16-1+1 DOWNTO 4*B_WIDTH/16+1) WHEN "0000000010000000",
      DOUT_REG_COMB1_9(6*B_WIDTH/16-1+1 DOWNTO 5*B_WIDTH/16+1) WHEN "0000000100000000",
      DOUT_REG_COMB1_9(7*B_WIDTH/16-1+1 DOWNTO 6*B_WIDTH/16+1) WHEN "0000001000000000",
      DOUT_REG_COMB1_9(8*B_WIDTH/16-1+1 DOWNTO 7*B_WIDTH/16+1) WHEN "0000010000000000",
      DOUT_REG_COMB1_9(9*B_WIDTH/16-1+1 DOWNTO 8*B_WIDTH/16+1) WHEN "0000100000000000",
      DOUT_REG_COMB1_9(10*B_WIDTH/16-1+1 DOWNTO 9*B_WIDTH/16+1) WHEN "0001000000000000",
      DOUT_REG_COMB1_9(11*B_WIDTH/16-1+1 DOWNTO 10*B_WIDTH/16+1) WHEN "0010000000000000",
      DOUT_REG_COMB1_9(12*B_WIDTH/16-1+1 DOWNTO 11*B_WIDTH/16+1) WHEN "0100000000000000",
      DOUT_REG_COMB1_9(13*B_WIDTH/16-1+1 DOWNTO 12*B_WIDTH/16+1) WHEN "1000000000000000",
      DOUT_REG_COMB1_9(14*B_WIDTH/16-1+1 DOWNTO 13*B_WIDTH/16+1) WHEN "0000000000000001",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB0_9 <=
      REG1_OUT WHEN "00000000000000001",
      REG0_OUT WHEN "00000000000000010",
      REG16_OUT WHEN "00000000000000100",
      REG15_OUT WHEN "00000000000001000",
      REG14_OUT WHEN "00000000000010000",
      REG13_OUT WHEN "00000000000100000",
      REG12_OUT WHEN "00000000001000000",
      REG11_OUT WHEN "00000000010000000",
      REG10_OUT WHEN "00000000100000000",
      REG9_OUT WHEN "00000001000000000",
      REG8_OUT WHEN "00000010000000000",
      REG7_OUT WHEN "00000100000000000",
      REG6_OUT WHEN "00001000000000000",
      REG5_OUT WHEN "00010000000000000",
      REG4_OUT WHEN "00100000000000000",
      REG3_OUT WHEN "01000000000000000",
      REG2_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB1_9 <=
      REG0_OUT WHEN "00000000000000001",
      REG16_OUT WHEN "00000000000000010",
      REG15_OUT WHEN "00000000000000100",
      REG14_OUT WHEN "00000000000001000",
      REG13_OUT WHEN "00000000000010000",
      REG12_OUT WHEN "00000000000100000",
      REG11_OUT WHEN "00000000001000000",
      REG10_OUT WHEN "00000000010000000",
      REG9_OUT WHEN "00000000100000000",
      REG8_OUT WHEN "00000001000000000",
      REG7_OUT WHEN "00000010000000000",
      REG6_OUT WHEN "00000100000000000",
      REG5_OUT WHEN "00001000000000000",
      REG4_OUT WHEN "00010000000000000",
      REG3_OUT WHEN "00100000000000000",
      REG2_OUT WHEN "01000000000000000",
      REG1_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 



    -- assignment for DOUT_10
    DOUT_10 <= DOUT_PART_10;
    WITH SEL_ADDR SELECT DOUT_PART_10 <=
      DOUT_REG_COMB0_10(3*B_WIDTH/16-1+1 DOWNTO 2*B_WIDTH/16+1) WHEN "0000000000000010",
      DOUT_REG_COMB0_10(4*B_WIDTH/16-1+1 DOWNTO 3*B_WIDTH/16+1) WHEN "0000000000000100",
      DOUT_REG_COMB0_10(5*B_WIDTH/16-1+1 DOWNTO 4*B_WIDTH/16+1) WHEN "0000000000001000",
      DOUT_REG_COMB0_10(6*B_WIDTH/16-1+1 DOWNTO 5*B_WIDTH/16+1) WHEN "0000000000010000",
      DOUT_REG_COMB0_10(7*B_WIDTH/16-1+1 DOWNTO 6*B_WIDTH/16+1) WHEN "0000000000100000",
      DOUT_REG_COMB0_10(8*B_WIDTH/16-1+1 DOWNTO 7*B_WIDTH/16+1) WHEN "0000000001000000",
      DOUT_REG_COMB0_10(9*B_WIDTH/16-1+1 DOWNTO 8*B_WIDTH/16+1) WHEN "0000000010000000",
      DOUT_REG_COMB0_10(10*B_WIDTH/16-1+1 DOWNTO 9*B_WIDTH/16+1) WHEN "0000000100000000",
      DOUT_REG_COMB0_10(11*B_WIDTH/16-1+1 DOWNTO 10*B_WIDTH/16+1) WHEN "0000001000000000",
      DOUT_REG_COMB0_10(12*B_WIDTH/16-1+1 DOWNTO 11*B_WIDTH/16+1) WHEN "0000010000000000",
      DOUT_REG_COMB0_10(13*B_WIDTH/16-1+1 DOWNTO 12*B_WIDTH/16+1) WHEN "0000100000000000",
      DOUT_REG_COMB0_10(14*B_WIDTH/16-1+1 DOWNTO 13*B_WIDTH/16+1) WHEN "0001000000000000",
      DOUT_REG_COMB0_10(15*B_WIDTH/16-1+1 DOWNTO 14*B_WIDTH/16+1) WHEN "0010000000000000",
      DOUT_REG_COMB1_10(0 DOWNTO 0) & DOUT_REG_COMB0_10(31 DOWNTO 15*B_WIDTH/16+1) WHEN "0100000000000000",
      DOUT_REG_COMB1_10(1*B_WIDTH/16-1+1 DOWNTO 0*B_WIDTH/16+1) WHEN "1000000000000000",
      DOUT_REG_COMB1_10(2*B_WIDTH/16-1+1 DOWNTO 1*B_WIDTH/16+1) WHEN "0000000000000001",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB0_10 <=
      REG12_OUT WHEN "00000000000000001",
      REG11_OUT WHEN "00000000000000010",
      REG10_OUT WHEN "00000000000000100",
      REG9_OUT WHEN "00000000000001000",
      REG8_OUT WHEN "00000000000010000",
      REG7_OUT WHEN "00000000000100000",
      REG6_OUT WHEN "00000000001000000",
      REG5_OUT WHEN "00000000010000000",
      REG4_OUT WHEN "00000000100000000",
      REG3_OUT WHEN "00000001000000000",
      REG2_OUT WHEN "00000010000000000",
      REG1_OUT WHEN "00000100000000000",
      REG0_OUT WHEN "00001000000000000",
      REG16_OUT WHEN "00010000000000000",
      REG15_OUT WHEN "00100000000000000",
      REG14_OUT WHEN "01000000000000000",
      REG13_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB1_10 <=
      REG11_OUT WHEN "00000000000000001",
      REG10_OUT WHEN "00000000000000010",
      REG9_OUT WHEN "00000000000000100",
      REG8_OUT WHEN "00000000000001000",
      REG7_OUT WHEN "00000000000010000",
      REG6_OUT WHEN "00000000000100000",
      REG5_OUT WHEN "00000000001000000",
      REG4_OUT WHEN "00000000010000000",
      REG3_OUT WHEN "00000000100000000",
      REG2_OUT WHEN "00000001000000000",
      REG1_OUT WHEN "00000010000000000",
      REG0_OUT WHEN "00000100000000000",
      REG16_OUT WHEN "00001000000000000",
      REG15_OUT WHEN "00010000000000000",
      REG14_OUT WHEN "00100000000000000",
      REG13_OUT WHEN "01000000000000000",
      REG12_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 



    -- assignment for DOUT_11
    DOUT_11 <= DOUT_PART_11;
    WITH SEL_ADDR SELECT DOUT_PART_11 <=
      DOUT_REG_COMB0_11(9*B_WIDTH/16-1+0 DOWNTO 8*B_WIDTH/16+0) WHEN "0000000000000010",
      DOUT_REG_COMB0_11(10*B_WIDTH/16-1+0 DOWNTO 9*B_WIDTH/16+0) WHEN "0000000000000100",
      DOUT_REG_COMB0_11(11*B_WIDTH/16-1+0 DOWNTO 10*B_WIDTH/16+0) WHEN "0000000000001000",
      DOUT_REG_COMB0_11(12*B_WIDTH/16-1+0 DOWNTO 11*B_WIDTH/16+0) WHEN "0000000000010000",
      DOUT_REG_COMB0_11(13*B_WIDTH/16-1+0 DOWNTO 12*B_WIDTH/16+0) WHEN "0000000000100000",
      DOUT_REG_COMB0_11(14*B_WIDTH/16-1+0 DOWNTO 13*B_WIDTH/16+0) WHEN "0000000001000000",
      DOUT_REG_COMB0_11(15*B_WIDTH/16-1+0 DOWNTO 14*B_WIDTH/16+0) WHEN "0000000010000000",
      DOUT_REG_COMB0_11(16*B_WIDTH/16-1+0 DOWNTO 15*B_WIDTH/16+0) WHEN "0000000100000000",
      DOUT_REG_COMB1_11(1*B_WIDTH/16-1+0 DOWNTO 0*B_WIDTH/16+0) WHEN "0000001000000000",
      DOUT_REG_COMB1_11(2*B_WIDTH/16-1+0 DOWNTO 1*B_WIDTH/16+0) WHEN "0000010000000000",
      DOUT_REG_COMB1_11(3*B_WIDTH/16-1+0 DOWNTO 2*B_WIDTH/16+0) WHEN "0000100000000000",
      DOUT_REG_COMB1_11(4*B_WIDTH/16-1+0 DOWNTO 3*B_WIDTH/16+0) WHEN "0001000000000000",
      DOUT_REG_COMB1_11(5*B_WIDTH/16-1+0 DOWNTO 4*B_WIDTH/16+0) WHEN "0010000000000000",
      DOUT_REG_COMB1_11(6*B_WIDTH/16-1+0 DOWNTO 5*B_WIDTH/16+0) WHEN "0100000000000000",
      DOUT_REG_COMB1_11(7*B_WIDTH/16-1+0 DOWNTO 6*B_WIDTH/16+0) WHEN "1000000000000000",
      DOUT_REG_COMB1_11(8*B_WIDTH/16-1+0 DOWNTO 7*B_WIDTH/16+0) WHEN "0000000000000001",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB0_11 <=
      REG7_OUT WHEN "00000000000000001",
      REG6_OUT WHEN "00000000000000010",
      REG5_OUT WHEN "00000000000000100",
      REG4_OUT WHEN "00000000000001000",
      REG3_OUT WHEN "00000000000010000",
      REG2_OUT WHEN "00000000000100000",
      REG1_OUT WHEN "00000000001000000",
      REG0_OUT WHEN "00000000010000000",
      REG16_OUT WHEN "00000000100000000",
      REG15_OUT WHEN "00000001000000000",
      REG14_OUT WHEN "00000010000000000",
      REG13_OUT WHEN "00000100000000000",
      REG12_OUT WHEN "00001000000000000",
      REG11_OUT WHEN "00010000000000000",
      REG10_OUT WHEN "00100000000000000",
      REG9_OUT WHEN "01000000000000000",
      REG8_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB1_11 <=
      REG6_OUT WHEN "00000000000000001",
      REG5_OUT WHEN "00000000000000010",
      REG4_OUT WHEN "00000000000000100",
      REG3_OUT WHEN "00000000000001000",
      REG2_OUT WHEN "00000000000010000",
      REG1_OUT WHEN "00000000000100000",
      REG0_OUT WHEN "00000000001000000",
      REG16_OUT WHEN "00000000010000000",
      REG15_OUT WHEN "00000000100000000",
      REG14_OUT WHEN "00000001000000000",
      REG13_OUT WHEN "00000010000000000",
      REG12_OUT WHEN "00000100000000000",
      REG11_OUT WHEN "00001000000000000",
      REG10_OUT WHEN "00010000000000000",
      REG9_OUT WHEN "00100000000000000",
      REG8_OUT WHEN "01000000000000000",
      REG7_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 



    -- assignment for DOUT_12
    DOUT_12 <= DOUT_PART_12;
    WITH SEL_ADDR SELECT DOUT_PART_12 <=
      DOUT_REG_COMB0_12(14*B_WIDTH/16-1+1 DOWNTO 13*B_WIDTH/16+1) WHEN "0000000000000010",
      DOUT_REG_COMB0_12(15*B_WIDTH/16-1+1 DOWNTO 14*B_WIDTH/16+1) WHEN "0000000000000100",
      DIN_IN(0 DOWNTO 0) & DOUT_REG_COMB0_12(31 DOWNTO 15*B_WIDTH/16+1) WHEN "0000000000001000",
      DOUT_REG_COMB1_12(1*B_WIDTH/16-1+1 DOWNTO 0*B_WIDTH/16+1) WHEN "0000000000010000",
      DOUT_REG_COMB1_12(2*B_WIDTH/16-1+1 DOWNTO 1*B_WIDTH/16+1) WHEN "0000000000100000",
      DOUT_REG_COMB1_12(3*B_WIDTH/16-1+1 DOWNTO 2*B_WIDTH/16+1) WHEN "0000000001000000",
      DOUT_REG_COMB1_12(4*B_WIDTH/16-1+1 DOWNTO 3*B_WIDTH/16+1) WHEN "0000000010000000",
      DOUT_REG_COMB1_12(5*B_WIDTH/16-1+1 DOWNTO 4*B_WIDTH/16+1) WHEN "0000000100000000",
      DOUT_REG_COMB1_12(6*B_WIDTH/16-1+1 DOWNTO 5*B_WIDTH/16+1) WHEN "0000001000000000",
      DOUT_REG_COMB1_12(7*B_WIDTH/16-1+1 DOWNTO 6*B_WIDTH/16+1) WHEN "0000010000000000",
      DOUT_REG_COMB1_12(8*B_WIDTH/16-1+1 DOWNTO 7*B_WIDTH/16+1) WHEN "0000100000000000",
      DOUT_REG_COMB1_12(9*B_WIDTH/16-1+1 DOWNTO 8*B_WIDTH/16+1) WHEN "0001000000000000",
      DOUT_REG_COMB1_12(10*B_WIDTH/16-1+1 DOWNTO 9*B_WIDTH/16+1) WHEN "0010000000000000",
      DOUT_REG_COMB1_12(11*B_WIDTH/16-1+1 DOWNTO 10*B_WIDTH/16+1) WHEN "0100000000000000",
      DOUT_REG_COMB1_12(12*B_WIDTH/16-1+1 DOWNTO 11*B_WIDTH/16+1) WHEN "1000000000000000",
      DOUT_REG_COMB1_12(13*B_WIDTH/16-1+1 DOWNTO 12*B_WIDTH/16+1) WHEN "0000000000000001",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB0_12 <=
      REG2_OUT WHEN "00000000000000001",
      REG1_OUT WHEN "00000000000000010",
      REG0_OUT WHEN "00000000000000100",
      REG16_OUT WHEN "00000000000001000",
      REG15_OUT WHEN "00000000000010000",
      REG14_OUT WHEN "00000000000100000",
      REG13_OUT WHEN "00000000001000000",
      REG12_OUT WHEN "00000000010000000",
      REG11_OUT WHEN "00000000100000000",
      REG10_OUT WHEN "00000001000000000",
      REG9_OUT WHEN "00000010000000000",
      REG8_OUT WHEN "00000100000000000",
      REG7_OUT WHEN "00001000000000000",
      REG6_OUT WHEN "00010000000000000",
      REG5_OUT WHEN "00100000000000000",
      REG4_OUT WHEN "01000000000000000",
      REG3_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB1_12 <=
      REG1_OUT WHEN "00000000000000001",
      REG0_OUT WHEN "00000000000000010",
      REG16_OUT WHEN "00000000000000100",
      REG15_OUT WHEN "00000000000001000",
      REG14_OUT WHEN "00000000000010000",
      REG13_OUT WHEN "00000000000100000",
      REG12_OUT WHEN "00000000001000000",
      REG11_OUT WHEN "00000000010000000",
      REG10_OUT WHEN "00000000100000000",
      REG9_OUT WHEN "00000001000000000",
      REG8_OUT WHEN "00000010000000000",
      REG7_OUT WHEN "00000100000000000",
      REG6_OUT WHEN "00001000000000000",
      REG5_OUT WHEN "00010000000000000",
      REG4_OUT WHEN "00100000000000000",
      REG3_OUT WHEN "01000000000000000",
      REG2_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 



    -- assignment for DOUT_13
    DOUT_13 <= DOUT_PART_13;
    WITH SEL_ADDR SELECT DOUT_PART_13 <=
      DOUT_REG_COMB0_13(2*B_WIDTH/16-1+1 DOWNTO 1*B_WIDTH/16+1) WHEN "0000000000000010",
      DOUT_REG_COMB0_13(3*B_WIDTH/16-1+1 DOWNTO 2*B_WIDTH/16+1) WHEN "0000000000000100",
      DOUT_REG_COMB0_13(4*B_WIDTH/16-1+1 DOWNTO 3*B_WIDTH/16+1) WHEN "0000000000001000",
      DOUT_REG_COMB0_13(5*B_WIDTH/16-1+1 DOWNTO 4*B_WIDTH/16+1) WHEN "0000000000010000",
      DOUT_REG_COMB0_13(6*B_WIDTH/16-1+1 DOWNTO 5*B_WIDTH/16+1) WHEN "0000000000100000",
      DOUT_REG_COMB0_13(7*B_WIDTH/16-1+1 DOWNTO 6*B_WIDTH/16+1) WHEN "0000000001000000",
      DOUT_REG_COMB0_13(8*B_WIDTH/16-1+1 DOWNTO 7*B_WIDTH/16+1) WHEN "0000000010000000",
      DOUT_REG_COMB0_13(9*B_WIDTH/16-1+1 DOWNTO 8*B_WIDTH/16+1) WHEN "0000000100000000",
      DOUT_REG_COMB0_13(10*B_WIDTH/16-1+1 DOWNTO 9*B_WIDTH/16+1) WHEN "0000001000000000",
      DOUT_REG_COMB0_13(11*B_WIDTH/16-1+1 DOWNTO 10*B_WIDTH/16+1) WHEN "0000010000000000",
      DOUT_REG_COMB0_13(12*B_WIDTH/16-1+1 DOWNTO 11*B_WIDTH/16+1) WHEN "0000100000000000",
      DOUT_REG_COMB0_13(13*B_WIDTH/16-1+1 DOWNTO 12*B_WIDTH/16+1) WHEN "0001000000000000",
      DOUT_REG_COMB0_13(14*B_WIDTH/16-1+1 DOWNTO 13*B_WIDTH/16+1) WHEN "0010000000000000",
      DOUT_REG_COMB0_13(15*B_WIDTH/16-1+1 DOWNTO 14*B_WIDTH/16+1) WHEN "0100000000000000",
      DOUT_REG_COMB1_13(0 DOWNTO 0) & DOUT_REG_COMB0_13(31 DOWNTO 15*B_WIDTH/16+1) WHEN "1000000000000000",
      DOUT_REG_COMB1_13(1*B_WIDTH/16-1+1 DOWNTO 0*B_WIDTH/16+1) WHEN "0000000000000001",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB0_13 <=
      REG13_OUT WHEN "00000000000000001",
      REG12_OUT WHEN "00000000000000010",
      REG11_OUT WHEN "00000000000000100",
      REG10_OUT WHEN "00000000000001000",
      REG9_OUT WHEN "00000000000010000",
      REG8_OUT WHEN "00000000000100000",
      REG7_OUT WHEN "00000000001000000",
      REG6_OUT WHEN "00000000010000000",
      REG5_OUT WHEN "00000000100000000",
      REG4_OUT WHEN "00000001000000000",
      REG3_OUT WHEN "00000010000000000",
      REG2_OUT WHEN "00000100000000000",
      REG1_OUT WHEN "00001000000000000",
      REG0_OUT WHEN "00010000000000000",
      REG16_OUT WHEN "00100000000000000",
      REG15_OUT WHEN "01000000000000000",
      REG14_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB1_13 <=
      REG12_OUT WHEN "00000000000000001",
      REG11_OUT WHEN "00000000000000010",
      REG10_OUT WHEN "00000000000000100",
      REG9_OUT WHEN "00000000000001000",
      REG8_OUT WHEN "00000000000010000",
      REG7_OUT WHEN "00000000000100000",
      REG6_OUT WHEN "00000000001000000",
      REG5_OUT WHEN "00000000010000000",
      REG4_OUT WHEN "00000000100000000",
      REG3_OUT WHEN "00000001000000000",
      REG2_OUT WHEN "00000010000000000",
      REG1_OUT WHEN "00000100000000000",
      REG0_OUT WHEN "00001000000000000",
      REG16_OUT WHEN "00010000000000000",
      REG15_OUT WHEN "00100000000000000",
      REG14_OUT WHEN "01000000000000000",
      REG13_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 



    -- assignment for DOUT_14
    DOUT_14 <= DOUT_PART_14;
    WITH SEL_ADDR SELECT DOUT_PART_14 <=
      DOUT_REG_COMB0_14(8*B_WIDTH/16-1+0 DOWNTO 7*B_WIDTH/16+0) WHEN "0000000000000010",
      DOUT_REG_COMB0_14(9*B_WIDTH/16-1+0 DOWNTO 8*B_WIDTH/16+0) WHEN "0000000000000100",
      DOUT_REG_COMB0_14(10*B_WIDTH/16-1+0 DOWNTO 9*B_WIDTH/16+0) WHEN "0000000000001000",
      DOUT_REG_COMB0_14(11*B_WIDTH/16-1+0 DOWNTO 10*B_WIDTH/16+0) WHEN "0000000000010000",
      DOUT_REG_COMB0_14(12*B_WIDTH/16-1+0 DOWNTO 11*B_WIDTH/16+0) WHEN "0000000000100000",
      DOUT_REG_COMB0_14(13*B_WIDTH/16-1+0 DOWNTO 12*B_WIDTH/16+0) WHEN "0000000001000000",
      DOUT_REG_COMB0_14(14*B_WIDTH/16-1+0 DOWNTO 13*B_WIDTH/16+0) WHEN "0000000010000000",
      DOUT_REG_COMB0_14(15*B_WIDTH/16-1+0 DOWNTO 14*B_WIDTH/16+0) WHEN "0000000100000000",
      DOUT_REG_COMB0_14(16*B_WIDTH/16-1+0 DOWNTO 15*B_WIDTH/16+0) WHEN "0000001000000000",
      DOUT_REG_COMB1_14(1*B_WIDTH/16-1+0 DOWNTO 0*B_WIDTH/16+0) WHEN "0000010000000000",
      DOUT_REG_COMB1_14(2*B_WIDTH/16-1+0 DOWNTO 1*B_WIDTH/16+0) WHEN "0000100000000000",
      DOUT_REG_COMB1_14(3*B_WIDTH/16-1+0 DOWNTO 2*B_WIDTH/16+0) WHEN "0001000000000000",
      DOUT_REG_COMB1_14(4*B_WIDTH/16-1+0 DOWNTO 3*B_WIDTH/16+0) WHEN "0010000000000000",
      DOUT_REG_COMB1_14(5*B_WIDTH/16-1+0 DOWNTO 4*B_WIDTH/16+0) WHEN "0100000000000000",
      DOUT_REG_COMB1_14(6*B_WIDTH/16-1+0 DOWNTO 5*B_WIDTH/16+0) WHEN "1000000000000000",
      DOUT_REG_COMB1_14(7*B_WIDTH/16-1+0 DOWNTO 6*B_WIDTH/16+0) WHEN "0000000000000001",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB0_14 <=
      REG8_OUT WHEN "00000000000000001",
      REG7_OUT WHEN "00000000000000010",
      REG6_OUT WHEN "00000000000000100",
      REG5_OUT WHEN "00000000000001000",
      REG4_OUT WHEN "00000000000010000",
      REG3_OUT WHEN "00000000000100000",
      REG2_OUT WHEN "00000000001000000",
      REG1_OUT WHEN "00000000010000000",
      REG0_OUT WHEN "00000000100000000",
      REG16_OUT WHEN "00000001000000000",
      REG15_OUT WHEN "00000010000000000",
      REG14_OUT WHEN "00000100000000000",
      REG13_OUT WHEN "00001000000000000",
      REG12_OUT WHEN "00010000000000000",
      REG11_OUT WHEN "00100000000000000",
      REG10_OUT WHEN "01000000000000000",
      REG9_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB1_14 <=
      REG7_OUT WHEN "00000000000000001",
      REG6_OUT WHEN "00000000000000010",
      REG5_OUT WHEN "00000000000000100",
      REG4_OUT WHEN "00000000000001000",
      REG3_OUT WHEN "00000000000010000",
      REG2_OUT WHEN "00000000000100000",
      REG1_OUT WHEN "00000000001000000",
      REG0_OUT WHEN "00000000010000000",
      REG16_OUT WHEN "00000000100000000",
      REG15_OUT WHEN "00000001000000000",
      REG14_OUT WHEN "00000010000000000",
      REG13_OUT WHEN "00000100000000000",
      REG12_OUT WHEN "00001000000000000",
      REG11_OUT WHEN "00010000000000000",
      REG10_OUT WHEN "00100000000000000",
      REG9_OUT WHEN "01000000000000000",
      REG8_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 



    -- assignment for DOUT_15
    DOUT_15 <= DOUT_PART_15;
    WITH SEL_ADDR SELECT DOUT_PART_15 <=
      DOUT_REG_COMB0_15(13*B_WIDTH/16-1+1 DOWNTO 12*B_WIDTH/16+1) WHEN "0000000000000010",
      DOUT_REG_COMB0_15(14*B_WIDTH/16-1+1 DOWNTO 13*B_WIDTH/16+1) WHEN "0000000000000100",
      DOUT_REG_COMB0_15(15*B_WIDTH/16-1+1 DOWNTO 14*B_WIDTH/16+1) WHEN "0000000000001000",
      DIN_IN(0 DOWNTO 0) & DOUT_REG_COMB0_15(31 DOWNTO 15*B_WIDTH/16+1) WHEN "0000000000010000",
      DOUT_REG_COMB1_15(1*B_WIDTH/16-1+1 DOWNTO 0*B_WIDTH/16+1) WHEN "0000000000100000",
      DOUT_REG_COMB1_15(2*B_WIDTH/16-1+1 DOWNTO 1*B_WIDTH/16+1) WHEN "0000000001000000",
      DOUT_REG_COMB1_15(3*B_WIDTH/16-1+1 DOWNTO 2*B_WIDTH/16+1) WHEN "0000000010000000",
      DOUT_REG_COMB1_15(4*B_WIDTH/16-1+1 DOWNTO 3*B_WIDTH/16+1) WHEN "0000000100000000",
      DOUT_REG_COMB1_15(5*B_WIDTH/16-1+1 DOWNTO 4*B_WIDTH/16+1) WHEN "0000001000000000",
      DOUT_REG_COMB1_15(6*B_WIDTH/16-1+1 DOWNTO 5*B_WIDTH/16+1) WHEN "0000010000000000",
      DOUT_REG_COMB1_15(7*B_WIDTH/16-1+1 DOWNTO 6*B_WIDTH/16+1) WHEN "0000100000000000",
      DOUT_REG_COMB1_15(8*B_WIDTH/16-1+1 DOWNTO 7*B_WIDTH/16+1) WHEN "0001000000000000",
      DOUT_REG_COMB1_15(9*B_WIDTH/16-1+1 DOWNTO 8*B_WIDTH/16+1) WHEN "0010000000000000",
      DOUT_REG_COMB1_15(10*B_WIDTH/16-1+1 DOWNTO 9*B_WIDTH/16+1) WHEN "0100000000000000",
      DOUT_REG_COMB1_15(11*B_WIDTH/16-1+1 DOWNTO 10*B_WIDTH/16+1) WHEN "1000000000000000",
      DOUT_REG_COMB1_15(12*B_WIDTH/16-1+1 DOWNTO 11*B_WIDTH/16+1) WHEN "0000000000000001",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB0_15 <=
      REG3_OUT WHEN "00000000000000001",
      REG2_OUT WHEN "00000000000000010",
      REG1_OUT WHEN "00000000000000100",
      REG0_OUT WHEN "00000000000001000",
      REG16_OUT WHEN "00000000000010000",
      REG15_OUT WHEN "00000000000100000",
      REG14_OUT WHEN "00000000001000000",
      REG13_OUT WHEN "00000000010000000",
      REG12_OUT WHEN "00000000100000000",
      REG11_OUT WHEN "00000001000000000",
      REG10_OUT WHEN "00000010000000000",
      REG9_OUT WHEN "00000100000000000",
      REG8_OUT WHEN "00001000000000000",
      REG7_OUT WHEN "00010000000000000",
      REG6_OUT WHEN "00100000000000000",
      REG5_OUT WHEN "01000000000000000",
      REG4_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 

    WITH SEL_REG_OUT SELECT DOUT_REG_COMB1_15 <=
      REG2_OUT WHEN "00000000000000001",
      REG1_OUT WHEN "00000000000000010",
      REG0_OUT WHEN "00000000000000100",
      REG16_OUT WHEN "00000000000001000",
      REG15_OUT WHEN "00000000000010000",
      REG14_OUT WHEN "00000000000100000",
      REG13_OUT WHEN "00000000001000000",
      REG12_OUT WHEN "00000000010000000",
      REG11_OUT WHEN "00000000100000000",
      REG10_OUT WHEN "00000001000000000",
      REG9_OUT WHEN "00000010000000000",
      REG8_OUT WHEN "00000100000000000",
      REG7_OUT WHEN "00001000000000000",
      REG6_OUT WHEN "00010000000000000",
      REG5_OUT WHEN "00100000000000000",
      REG4_OUT WHEN "01000000000000000",
      REG3_OUT WHEN "10000000000000000",
      (OTHERS => '0') WHEN OTHERS; 



    -- selection of the correct registers to create output   
    SELECTION_REG : PROCESS(CLK)
    BEGIN
        IF RISING_EDGE(CLK) THEN
            IF RESET = '1' THEN
                SEL_REG_OUT <= "10000000000000000";
            ELSE
                IF SEL_ADDR = "0000000000000001" AND CNT_DONE_INIT = '1' THEN
                    SEL_REG_OUT <= SEL_REG_OUT(15 DOWNTO 0) & SEL_REG_OUT(16);
                ELSE 
                    SEL_REG_OUT <= SEL_REG_OUT;
                END IF;
            END IF;
        END IF;
    END PROCESS;
    ------------------------------------------------------------------------------
  

    -- REGISTER ------------------------------------------------------------------
    -- generate selection signal to read from lower or upper part of the polynomial    
    SELECTION_ADDR : PROCESS(CLK)
    BEGIN
        IF RISING_EDGE(CLK) THEN
            IF RESET = '1' THEN
                SEL_ADDR <= "0000000000000001";
            ELSE
                IF SEL_ADDR_EN = '1' THEN
                    SEL_ADDR <= SEL_ADDR(14 DOWNTO 0) & SEL_ADDR(15);
                ELSE 
                    SEL_ADDR <= SEL_ADDR;
                END IF;
            END IF;
        END IF;
    END PROCESS;
    
    -- select the correct part of the polynomial
    WITH SEL_ADDR SELECT ADDR_IN <=
      CNT_OUT_0 WHEN "0000000000000001",
      CNT_OUT_1 WHEN "0000000000000010",
      CNT_OUT_2 WHEN "0000000000000100",
      CNT_OUT_3 WHEN "0000000000001000",
      CNT_OUT_4 WHEN "0000000000010000",
      CNT_OUT_5 WHEN "0000000000100000",
      CNT_OUT_6 WHEN "0000000001000000",
      CNT_OUT_7 WHEN "0000000010000000",
      CNT_OUT_8 WHEN "0000000100000000",
      CNT_OUT_9 WHEN "0000001000000000",
      CNT_OUT_10 WHEN "0000010000000000",
      CNT_OUT_11 WHEN "0000100000000000",
      CNT_OUT_12 WHEN "0001000000000000",
      CNT_OUT_13 WHEN "0010000000000000",
      CNT_OUT_14 WHEN "0100000000000000",
      CNT_OUT_15 WHEN "1000000000000000",
      (OTHERS => '0') WHEN OTHERS;

    -- registers to hold previous read words   
    SELECTION_REG_EN : PROCESS(CLK)
    BEGIN
        IF RISING_EDGE(CLK) THEN
            IF RESET = '1' THEN
                REG_EN <= "00000000000000001";
            ELSE
                IF SEL_REG_EN = '1' THEN
                    REG_EN <= REG_EN(15 DOWNTO 0) & REG_EN(16);
                ELSE 
                    REG_EN <= REG_EN;
                END IF;
            END IF;
        END IF;
    END PROCESS;
      
    REG_IN  <= DIN_IN;
  
    REG0 : ENTITY work.RegisterFDRE GENERIC MAP (SIZE => B_WIDTH)
    PORT MAP(D => REG_IN, Q => REG0_OUT, CLK => CLK, EN => REG_EN(0), RST => RESET);
    REG1 : ENTITY work.RegisterFDRE GENERIC MAP (SIZE => B_WIDTH)
    PORT MAP(D => REG_IN, Q => REG1_OUT, CLK => CLK, EN => REG_EN(1), RST => RESET);
    REG2 : ENTITY work.RegisterFDRE GENERIC MAP (SIZE => B_WIDTH)
    PORT MAP(D => REG_IN, Q => REG2_OUT, CLK => CLK, EN => REG_EN(2), RST => RESET);
    REG3 : ENTITY work.RegisterFDRE GENERIC MAP (SIZE => B_WIDTH)
    PORT MAP(D => REG_IN, Q => REG3_OUT, CLK => CLK, EN => REG_EN(3), RST => RESET);
    REG4 : ENTITY work.RegisterFDRE GENERIC MAP (SIZE => B_WIDTH)
    PORT MAP(D => REG_IN, Q => REG4_OUT, CLK => CLK, EN => REG_EN(4), RST => RESET);
    REG5 : ENTITY work.RegisterFDRE GENERIC MAP (SIZE => B_WIDTH)
    PORT MAP(D => REG_IN, Q => REG5_OUT, CLK => CLK, EN => REG_EN(5), RST => RESET);
    REG6 : ENTITY work.RegisterFDRE GENERIC MAP (SIZE => B_WIDTH)
    PORT MAP(D => REG_IN, Q => REG6_OUT, CLK => CLK, EN => REG_EN(6), RST => RESET);
    REG7 : ENTITY work.RegisterFDRE GENERIC MAP (SIZE => B_WIDTH)
    PORT MAP(D => REG_IN, Q => REG7_OUT, CLK => CLK, EN => REG_EN(7), RST => RESET);
    REG8 : ENTITY work.RegisterFDRE GENERIC MAP (SIZE => B_WIDTH)
    PORT MAP(D => REG_IN, Q => REG8_OUT, CLK => CLK, EN => REG_EN(8), RST => RESET);
    REG9 : ENTITY work.RegisterFDRE GENERIC MAP (SIZE => B_WIDTH)
    PORT MAP(D => REG_IN, Q => REG9_OUT, CLK => CLK, EN => REG_EN(9), RST => RESET);
    REG10 : ENTITY work.RegisterFDRE GENERIC MAP (SIZE => B_WIDTH)
    PORT MAP(D => REG_IN, Q => REG10_OUT, CLK => CLK, EN => REG_EN(10), RST => RESET);
    REG11 : ENTITY work.RegisterFDRE GENERIC MAP (SIZE => B_WIDTH)
    PORT MAP(D => REG_IN, Q => REG11_OUT, CLK => CLK, EN => REG_EN(11), RST => RESET);
    REG12 : ENTITY work.RegisterFDRE GENERIC MAP (SIZE => B_WIDTH)
    PORT MAP(D => REG_IN, Q => REG12_OUT, CLK => CLK, EN => REG_EN(12), RST => RESET);
    REG13 : ENTITY work.RegisterFDRE GENERIC MAP (SIZE => B_WIDTH)
    PORT MAP(D => REG_IN, Q => REG13_OUT, CLK => CLK, EN => REG_EN(13), RST => RESET);
    REG14 : ENTITY work.RegisterFDRE GENERIC MAP (SIZE => B_WIDTH)
    PORT MAP(D => REG_IN, Q => REG14_OUT, CLK => CLK, EN => REG_EN(14), RST => RESET);
    REG15 : ENTITY work.RegisterFDRE GENERIC MAP (SIZE => B_WIDTH)
    PORT MAP(D => REG_IN, Q => REG15_OUT, CLK => CLK, EN => REG_EN(15), RST => RESET);
    REG16 : ENTITY work.RegisterFDRE GENERIC MAP (SIZE => B_WIDTH)
    PORT MAP(D => REG_IN, Q => REG16_OUT, CLK => CLK, EN => REG_EN(16), RST => RESET);
    ------------------------------------------------------------------------------

    -- FSM -----------------------------------------------------------------------
    FSM : PROCESS(CLK)
    BEGIN
        IF RISING_EDGE(CLK) THEN
            CASE STATE IS
                
                ----------------------------------------------
                WHEN S_RESET        =>
                    -- GLOBAL ----------
                    DONE                    <= '0';
                
                    -- COUNTER ---------
                    CNT_EN_OUT              <= '0';
                    CNT_RST_OUT             <= '1';
                    
                    CNT_EN_INIT             <= '0';
                    CNT_RST_INIT            <= '1';
                    
                    CNT_RST                 <= '1';
                    
                    -- CONTROL ---------
                    SEL_REG_EN              <= '0';
                    SEL_ADDR_EN             <= '0'; 
                    
                    -- BRAM ------------
                    REN_IN                  <= '0';
                    WEN_OUT                 <= '0';
                    
                    -- TRANSITION ------
                    IF (ENABLE = '1') THEN                      
                        STATE               <= S_INIT0;
                    ELSE
                        STATE               <= S_RESET;
                    END IF;
                ----------------------------------------------

                ----------------------------------------------
                WHEN S_INIT0  =>
                    -- GLOBAL ----------
                    DONE                    <= '0';
                
                    -- COUNTER ---------
                    CNT_EN_OUT              <= '0';
                    CNT_RST_OUT             <= '1';

                    CNT_EN_INIT             <= '1';
                    CNT_RST_INIT            <= '0';
                                        
                    CNT_RST                 <= '0';
                    
                    -- CONTROL ---------
                    SEL_REG_EN              <= '0';
                    SEL_ADDR_EN             <= '1';                
                    
                    -- BRAM ------------
                    REN_IN                  <= '1';
                    WEN_OUT                 <= '0';
                                      
                    -- TRANSITION ------
                    STATE                   <= S_INIT1;
                ----------------------------------------------    

                ----------------------------------------------
                WHEN S_INIT1  =>
                    -- GLOBAL ----------
                    DONE                    <= '0';
                
                    -- COUNTER ---------
                    CNT_EN_OUT              <= '0';
                    CNT_RST_OUT             <= '1';
                    
                    CNT_EN_INIT             <= '1';
                    CNT_RST_INIT            <= '0';
                    
                    CNT_RST                 <= '0';
                    
                    -- CONTROL ---------
                    SEL_REG_EN              <= '1';
                    SEL_ADDR_EN             <= '1';                
                    
                    -- BRAM ------------
                    REN_IN                  <= '1';
                    WEN_OUT                 <= '0';
                                      
                    -- TRANSITION ------
                    --STATE <= S_INIT2;
                    IF (CNT_DONE_INIT = '1') THEN
                        STATE               <= S_WRITE;
                    ELSE
                        STATE               <= S_INIT1;
                    END IF;
                ----------------------------------------------
                                
                ----------------------------------------------
                WHEN S_WRITE  =>
                    -- GLOBAL ----------
                    DONE                    <= '0';
                
                    -- COUNTER ---------
                    CNT_EN_OUT              <= '1';
                    CNT_RST_OUT             <= '0';
                    
                    CNT_EN_INIT             <= '0';
                    CNT_RST_INIT            <= '0';
                    
                    CNT_RST                 <= '0';
                    
                    -- CONTROL ---------
                    SEL_REG_EN              <= '1';
                    SEL_ADDR_EN             <= '1';                
                    
                    -- BRAM ------------
                    REN_IN                  <= '1';
                    WEN_OUT                 <= '1';   
                                                        
                    -- TRANSITION ------
                    IF (CNT_DONE_OUT = '1') THEN
                        STATE               <= S_DONE;
                    ELSE
                        STATE               <= S_WRITE;
                    END IF;
                ---------------------------------------------- 
                                                                
                ----------------------------------------------
                WHEN S_DONE         =>
                    -- GLOBAL ----------
                    DONE                    <= '1';
                
                    -- COUNTER ---------
                    CNT_EN_OUT              <= '0';
                    CNT_RST_OUT             <= '1';

                    
                    CNT_EN_INIT             <= '0';
                    CNT_RST_INIT            <= '1';
                                        
                    CNT_RST                 <= '1';
                    
                    -- CONTROL ---------
                    SEL_REG_EN              <= '0';
                    SEL_ADDR_EN             <= '0';                
                    
                    -- BRAM ------------
                    REN_IN                  <= '0';
                    WEN_OUT                 <= '0';
                                        
                    -- TRANSITION ------
                    STATE                   <= S_RESET;
                ----------------------------------------------
                                
            END CASE;
        END IF;
    END PROCESS;    
    ------------------------------------------------------------------------------

END Behavioral;
